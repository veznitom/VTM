package global_variables is
	constant XLEN : integer := 32;
end package global_variables;