module Loader (
  input wire [31:0][2] instr_in,
  input wire stop,
  output reg [31:0][2] instr_out,
  output reg ready
);

endmodule
