module reorder_buffer #(
    parameter int XLEN = 32
) (
    global_signals_if gsi,
    pc_interface_if pc,
    common_data_bus_if cdb[2],
    instr_issue_if iii[2]
);
    TODO();
endmodule
