module branch #(
    parameter int XLEN = 32
) (
    station_unit_if exec_feed,

    output logic [XLEN-1:0] store_result, jump_result
);
    TODO();
endmodule
