module cache #(
    parameter int XLEN = 32
) (
    global_signals_if gsi,

    cache_bus_if cache_bus,
    cache_memory_bus_if memory_bus,
    common_data_bus_if cdb[2]
);
    TODO();
endmodule
