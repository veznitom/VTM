package flags
  typedef logic [7:0] flag;

 const flag REG_WRITE = 8'b00000001;
 const flag CACHE_WRITE = 8'b00000001;
endpackage