module register_file #(
    parameter int XLEN = 32
) (
    global_signals_if gsi,
    register_query_if queries[2],
    register_values_if reg_reses[2]
);
    TODO();
endmodule
