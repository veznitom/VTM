module ip_renamer (
    input clock,
    input reset
);

endmodule
