// Copyright (c) 2024 veznitom

`default_nettype none
import pkg_defines::*;
module RenameManager (
  IntfCSB.notag cs,

  input  wire       i_get,
  output wire [5:0] o_rnn,
  output wire [1:0] o_left
);
endmodule
