module data_cache #(
    parameter int XLEN = 32
) (
    global_signals_if gsi,

    data_cache_bus_if data_bus,
    data_memory_bus_if mem_bus,

    common_data_bus_if cdb[2]
);
    TODO();
endmodule
