package global_variables;
  integer XLEN = 32;
endpackage : global_variables
