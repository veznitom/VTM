package global_variables;
  localparam integer XLEN = 32;
endpackage : global_variables
