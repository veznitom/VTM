module cache #(
    parameter int XLEN = 32
) (
    global_signals_if gsi,

    cache_bus_if cache_bus,
    data_memory_bus_if mem_bus,

    common_data_bus_if cdb[2]
);
    TODO();
endmodule
