module load_store #(
    parameter int XLEN = 32
) (
    station_unit_if exec_feed,
    data_cache_bus_if data_bus,

    output logic [XLEN-1:0] result
);
    TODO();
endmodule
