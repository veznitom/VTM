// Copyright (c) 2024 veznitom

`default_nettype none
import pkg_defines::*;
module Control (
  input wire i_clock,
  input wire i_reset
);

endmodule
