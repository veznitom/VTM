module register_file #(
    parameter int XLEN = 32
) (
    global_signals_if gsi,
    register_query_if query[2],
    register_values_if reg_val[2],
    debug_interface_if debug
);
    TODO();
endmodule
