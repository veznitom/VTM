package vtm_enums is
  type INSTR_NAME_E is (TMP);
  type INSTR_TYPE_E is (AL);
end package vtm_enums;

package vtm_records is

end package vtm_records;
