module program_counter #(
    parameter int XLEN = 32
) (
    pc_interface_if inter
);
  TODO();
endmodule
