module mem_mng_unit (
    global_signals_if gsi,
    data_memory_bus_if data_bus,
    instr_memory_bus_if instr_bus,
    memory_bus_if memory_bus
);
    TODO();
endmodule
