module ip_control (
    input clock,
    input reset
);

endmodule
