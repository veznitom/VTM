module pc (
    pc_interface_if inter
);
    TODO();
endmodule
